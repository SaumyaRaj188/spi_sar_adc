/*
 * Module: adc_spi_slave
 * Description: SPI Slave Interface matching the README.md register map.
 * Handles Register R/W, EOC latching, and status updates.
 */
module adc_spi_slave (
    // System Interface
    input           clk,            // System Clock
    input           reset_,         // Active-low Reset

    // SPI Interface
    input           cs,             // Chip Select
    input           sck,            // SPI Clock
    input           mosi,           // Master Out Slave In
    output          miso,           // Master In Slave Out

    // Hardware Interface (Connections to Top Level/ADC)
    input  [11:0]   adc_data_in,    // Live Data from ADC
    input           adc_busy_in,    // Live Busy Status from ADC
    input           adc_eoc_pulse,  // Pulse from ADC when conversion finishes (Sets EOC)
    input           hw_clear_start, // Signal from Top Level to clear the START bit
    output [11:0]   ctrl_reg_out,   // Expose Control Register to Top Level
    output          eoc_flag_out    // Expose EOC status for Interrupts
);

    // -- Address Map --
    localparam ADDR_CTRL   = 2'b00;
    localparam ADDR_STATUS = 2'b01;
    localparam ADDR_DATA   = 2'b10;
    localparam ADDR_INFO   = 2'b11;

    // -- Command Map --
    localparam CMD_READ  = 2'b00;
    localparam CMD_WRITE = 2'b01;
    localparam CMD_SET   = 2'b10;
    localparam CMD_CLEAR = 2'b11;

    // -- Internal Registers --
    reg [11:0] ctrl_reg;     
    reg        eoc_latch;    
    reg [11:0] data_reg;     
    reg [11:0] info_reg;     

    // -- SPI Logic Signals --
    reg [1:0]  state;
    reg [4:0]  bit_cnt;
    reg [15:0] shift_reg;
    reg [11:0] miso_buffer;
    
    // SCK Synchronization
    reg sck_s1, sck_s2;
    wire sck_rise;
    wire sck_fall;

    assign sck_rise = (sck_s1 && !sck_s2);
    assign sck_fall = (!sck_s1 && sck_s2);

    // Frame Parsing
    wire [1:0]  cmd;
    wire [1:0]  addr;
    wire [11:0] pay;
    
    assign cmd  = shift_reg[15:14];
    assign addr = shift_reg[13:12];
    assign pay  = shift_reg[11:0];

    // -- State Machine --
    localparam S_IDLE  = 2'b00;
    localparam S_SHIFT = 2'b01;
    localparam S_LATCH = 2'b10;

    // -- Assignments --
    assign ctrl_reg_out = ctrl_reg;
    assign eoc_flag_out = eoc_latch; 
    assign miso         = cs ? 1'bz : miso_buffer[11];

    // -- SCK Synchronizer --
    always @(posedge clk or negedge reset_) begin
        if(!reset_) begin
            sck_s1 <= 0; sck_s2 <= 0;
        end else begin
            sck_s1 <= sck; sck_s2 <= sck_s1;
        end
    end

    // -- Main State Machine & Datapath --
    always @(posedge clk or negedge reset_) begin
        if(!reset_) begin
            state       <= S_IDLE;
            ctrl_reg    <= 12'h0;
            data_reg    <= 12'h0;
            info_reg    <= 12'h00A; 
            eoc_latch   <= 1'b0;
            bit_cnt     <= 0;
            shift_reg   <= 0;
            miso_buffer <= 0;
        end else begin
            
            // 1. EOC Management
            if (adc_eoc_pulse) begin
                eoc_latch <= 1'b1;
            end
            
            // 2. Hardware Clear of START bit
            if (hw_clear_start) begin
                ctrl_reg[1] <= 1'b0; 
            end

            case(state)
                S_IDLE: begin
                    bit_cnt <= 0;
                    data_reg <= adc_data_in; // Update Live Data
                    if(!cs) state <= S_SHIFT;
                end

                S_SHIFT: begin
                    // Priority Check: CS de-assertion terminates frame
                    if(cs) begin
                         // OPTIONAL: If we have exactly 16 bits when CS goes high, we could latch.
                         // But for Mode 0, we usually latch on the last clock edge.
                         // For safety, we just go to IDLE here.
                         state <= S_IDLE; 
                    end else if(sck_rise) begin
                        // Shift In
                        shift_reg <= {shift_reg[14:0], mosi}; 
                        bit_cnt   <= bit_cnt + 1;
                        
                        // FIX: Transition to LATCH on the 16th edge (when count is 15 -> 16)
                        if (bit_cnt == 15) begin
                            state <= S_LATCH;
                        end
                    end

                    // Shift Out (MISO) on Falling Edge
                    if(!cs && sck_fall) begin
                         miso_buffer <= {miso_buffer[10:0], 1'b0};
                    end

                    // Pre-load MISO buffer logic (after 4 bits)
                    // We look at bit_cnt == 4 because we just incremented it on rise.
                    // But we need to load it before the next fall shift.
                    if(!cs && bit_cnt == 4 && sck_fall) begin 
                         // Note: We access shift_reg directly. The 4 bits are at [3:0] of shift_reg
                         // because we shift left. Wait, shift_reg shifts in at LSB.
                         // After 4 shifts: [15:4] is old garbage, [3:0] is the new CMD/ADDR.
                         // Wait, code says `cmd = shift_reg[15:14]`. That implies shift_reg holds result at END.
                         // During shift, the bits are moving.
                         // Let's rely on the previous logic which worked for Read.
                         // Actually, simpler logic: Only load MISO buffer if we are doing a read.
                         // The previous logic was slightly fragile regarding shift position.
                         
                         // Simplified MISO Load:
                         // We can't easily parse CMD/ADDR mid-stream without complex indexing.
                         // For this fix, I will focus on the WRITE functionality working first.
                         // The READ functionality relies on fully received bits.
                         
                         // Let's stick to the previous working MISO logic, just adjusted:
                         if (shift_reg[3:2] == CMD_READ) begin 
                           case(shift_reg[1:0])
                                ADDR_CTRL:   miso_buffer <= ctrl_reg;
                                ADDR_STATUS: miso_buffer <= {10'b0, adc_busy_in, eoc_latch};
                                ADDR_DATA:   miso_buffer <= data_reg;
                                ADDR_INFO:   miso_buffer <= info_reg;
                           endcase
                        end
                    end
                end

                S_LATCH: begin
                    // We arrived here because we received 16 bits.
                    state <= S_IDLE; 
                    
                    // Execute Write Commands
                    // Note: The shift_reg is now fully populated.
                    if (addr == ADDR_CTRL) begin
                        case(cmd)
                            CMD_WRITE: ctrl_reg <= pay;
                            CMD_SET:   ctrl_reg <= ctrl_reg | pay;
                            CMD_CLEAR: ctrl_reg <= ctrl_reg & ~pay;
                        endcase
                    end
                    
                    if (cmd == CMD_READ && addr == ADDR_STATUS) begin
                        eoc_latch <= 1'b0;
                    end
                end
            endcase
        end
    end

endmodule